// MatrixDisplay.sv
// Output signals to the Matrix display
// Bryce Adam
// Mar 05, 2024